`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name:    pillar_con 
// Description: 
//////////////////////////////////////////////////////////////////////////////////
module pillar_con(input reg [2:0]stage, 
						input reg [6:0]speed, 
						output reg [9:0]pillar_x, 
						output reg [8:0]pillar_y
    );


endmodule
